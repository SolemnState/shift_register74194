`timescale 1ns / 1ps
//  SPB SUAI
//Group 1641
// Authors:   Filippov K. and Denisov D. 
// XOR module with 2 inputs and 1 output.
module XOR(
    input a,
    input b,
    output c
    );
    assign c=a^b;
endmodule
